----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/02/2022 05:14:41 PM
-- Design Name: 
-- Module Name: load - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity load is
  Port (b : IN std_logic_vector(7 downto 0); c : IN std_logic; S : OUT std_logic_vector(8 downto 0));
end load;

architecture Behavioral of load is

Signal beta : std_logic_vector(7 downto 0);

begin
beta<=b;
S<=c&beta;



end Behavioral;
